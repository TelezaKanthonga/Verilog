module hello;

initial
begin
  $display("Hello World \n\n");
end

endmodule
